/********************************************************
** Pulse Average Blocks: 200-223
********************************************************/
localparam [7:0] SR_PULSE_LENGTH = 200;
localparam [7:0] SR_PULSE_NUM_AVG = 201;

/* Control readback registers */
localparam [7:0] RB_PULSE_LENGTH         = 0;
